/*
Assignment 5
Problem no: 3
Semester: 5th
Group: 28
Members: 
Aryan Singh (19CS30007)
Abhinandan De (19CS10069)
*/

`timescale 1ns/1ns

`ifndef _UnsignedCmp_v_
`define _UnsignedCmp_v_
`include "Dff.v"

// module dff_struct(D, Clk, Reset, Q);

module UnsignedCmp(
        input reset,

        input clk,
        output reg res
    );
    
    wire ;

endmodule

`endif 
